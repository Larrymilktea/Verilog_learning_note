//=======================================================
//  通用波形測試模板 (for Icarus Verilog + GTKWave)
//=======================================================

`timescale 1ns/1ps

module tb;           // tb = testbench (頂層模組)
  reg clk;           // 宣告時脈
  reg rst;           // 宣告 reset 訊號
  reg a, b;          // 測試輸入
  wire y;            // 被測模組輸出

  //=======================================================
  // 例化（instantiation）— 你要測的模組
  //=======================================================
  and_gate uut (
    .a(a),
    .b(b),
    .y(y)
  );

  //=======================================================
  // 產生波形輸出 (必要的兩行)
  //=======================================================
  initial begin
    $dumpfile("test.vcd");    // 指定輸出波形檔案
    $dumpvars(0, tb);         // 把 tb 模組的所有信號都記錄下來
  end

  //=======================================================
  // 產生時脈與測試輸入
  //=======================================================
  initial begin
    clk = 0; rst = 1; a = 0; b = 0;
    #5  rst = 0;
    #10 a = 1; b = 0;
    #10 a = 0; b = 1;
    #10 a = 1; b = 1;
    #10 $finish;
  end

  always #5 clk = ~clk;  // 10ns 時脈週期
endmodule


//=======================================================
//  被測模組 (例: AND Gate)
//=======================================================
module and_gate(input a, input b, output y);
  assign y = a & b;
endmodule
